

module task_2(
	input a, b, c, d,
    output q );

assign q = c | b;

endmodule